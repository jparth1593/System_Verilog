
//typedef class fa_intf;

class fa_cfg;

static mailbox gentobfm = new();

static virtual fa_intf svif;  // declaration of interface

endclass