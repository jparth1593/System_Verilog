interface fa_intf;
// define port name as per fa_tx
	logic  a;
	logic  b;
	logic  cin;
	logic  s;
	logic  c_out;

endinterface